module ram_fibx(A,Rd,Wd,Wen);
    input [15:0] A;
    input [15:0] Wd;
    output [15:0] Rd;
    

    if (Wen)



16'hD900
16'hD907
16'h2501
16'h2500
16'h60C0
16'h8030
16'h0683
16'h2430
16'hAC14
16'h70C0
16'h94C0
16'h1B00


endmodule
